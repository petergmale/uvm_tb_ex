
package env_pkg;

endpackage : env_pkg
