
package vseq_lib_pkg;

endpackage : vseq_lib_pkg
