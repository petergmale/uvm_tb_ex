
package seq_lib_pkg;

endpackage : seq_lib_pkg
