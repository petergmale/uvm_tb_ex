

module DUT (
        input   clk,
        input   rstn,
        input   sig1,
        input   sig2,
        output  sig3
    );

endmodule

