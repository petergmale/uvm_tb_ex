
interface a_if( input clk, rstn);

  logic   sig1;
  logic   sig2;
  logic   sig3;



  //- Protocol Assertions
    
endinterface


