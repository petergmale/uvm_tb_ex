
package agent_pkg;

endpackage : agent_pkg
